library ieee;
use ieee.std_logic_1164.all;

entity uart is 

    
end entity;

architecture logic of uart is 
begin

end architecture;