library ieee;
use ieee.std_logic_1164.all;

entity led_driver is 

end entity;

architecture logic of led_driver is 
begin

end architecture;