library ieee;
use ieee.std_logic_1164.all;

entity edge_divider is 

end entity;

architecture logic of edge_divider is 
begin


end architecture;