library ieee;
use ieee.std_logic_1164.all;

entity blinky is 

end entity;

architecture logic of blinky is 
begin 

end architecture;